library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use STD.TEXTIO.ALL;
use IEEE.STD_LOGIC_TEXTIO.ALL;

entity one_shot_tb is
end one_shot_tb;

architecture behav of one_shot_tb is
	component one_shot
        Port (
	sys_clk, reset, trigger_i    : in  STD_LOGIC;
	pulse_o    : out STD_LOGIC);
	end component;
    
	signal sys_clk, reset, trigger_i   : STD_LOGIC := '0';
	signal pulse_o   : STD_LOGIC;
    
	constant clk_period : time := 20 ns;
	file output_file : text;
    
begin
	uut: one_shot
	Port map (
	sys_clk   => sys_clk,
	reset     => reset,
	trigger_i => trigger_i,
	pulse_o   => pulse_o);
    
clk_process: process
begin
	sys_clk <= '0';
        wait for clk_period/2;
        sys_clk <= '1';
        wait for clk_period/2;
end process;

file_write: process(sys_clk)
	variable file_line : line;
	variable file_status : file_open_status;
	variable first_edge : boolean := true;
begin
	if rising_edge(sys_clk) then
		if first_edge then
                file_open(file_status, output_file, "one_shot_results.csv", write_mode);
                write(file_line, string'("Time_ns,Reset,Trigger_i,Pulse_o"));
                writeline(output_file, file_line);
                first_edge := false;
            	end if;
            
	write(file_line, integer'image(now / 1 ns));
	write(file_line, string'(","));
	write(file_line, std_logic'image(reset));
	write(file_line, string'(","));
	write(file_line, std_logic'image(trigger_i));
	write(file_line, string'(","));
	write(file_line, std_logic'image(pulse_o));
	writeline(output_file, file_line);
        end if;
end process;

bench_process: process
begin
        report "=== Starting One-Shot Testbench ===" severity note;
        reset <= '1';
        trigger_i <= '0';
        wait for 100 ns;
        report "Test 1: Reset applied" severity note;
        
        reset <= '0';
        wait for 50 ns;
        report "Test 1: Reset released" severity note;
        
        report "Test 2: Short trigger pulse (30 ns)" severity note;
        trigger_i <= '1';
        wait for 30 ns;
        trigger_i <= '0';
        wait for 100 ns;
        report "Test 2: Pulse_o = " & std_logic'image(pulse_o) severity note;
        
        report "Test 3: Long trigger pulse (200 ns)" severity note;
        trigger_i <= '1';
        wait for 200 ns;
        trigger_i <= '0';
        wait for 100 ns;
        report "Test 3: Pulse_o = " & std_logic'image(pulse_o) severity note;
        
        report "Test 4: Multiple trigger pulses" severity note;
        trigger_i <= '1';
        wait for 50 ns;
        trigger_i <= '0';
        wait for 80 ns;
        
        trigger_i <= '1';
        wait for 40 ns;
        trigger_i <= '0';
        wait for 100 ns;
        report "Test 4: Multiple pulses completed" severity note;
        
        file_close(output_file);
        report "=== Simulation Complete. Data saved to one_shot_results.csv ===" severity note;
        wait;
end process;
    
end behav;