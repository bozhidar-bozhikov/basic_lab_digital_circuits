library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity one_shot is
    Port (
        sys_clk, reset, trigger_i    : in  STD_LOGIC;
        pulse_o    : out STD_LOGIC
    );
end one_shot;

architecture behav of one_shot is
    signal state, next_state      : std_logic := '0';
    
begin
    state_memory: process(reset, sys_clk)
    begin
        if reset = '1' then
            state <= '0';
        elsif rising_edge(sys_clk) then
            state <= next_state;
        end if;
    end process state_memory;
    
    next_state_process: process(reset, trigger_i, state)
    begin
        if reset = '1' then
            next_state <= '0';
        elsif rising_edge(trigger_i) then
            next_state <= '1';
        elsif state = '1' then
            next_state <= '0';
        else
            next_state <= state;
        end if;
    end process next_state_process;
    
    pulse_o <= state;
    
end behav;